`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369A - Computer Architecture
// Laboratory 
// Module - InstructionMemory_tb.v
// Description - Test the 'InstructionMemory_tb.v' module.
////////////////////////////////////////////////////////////////////////////////

module InstructionMemory_tb(); 

    wire [31:0] Instruction;

    reg [31:0] Address;

	InstructionMemory u0(
		.Address(Address),
        .Instruction(Instruction)
	);

	initial begin
	
    	/* Please fill in the implementation here... */
		Address = 32'h00000001;
    		#10; 
    		Address = 32'h00000002;
    		#10; 
    		Address = 32'h00000003;
    		#10; 
    		Address = 32'h00000004;
    		#10; 
    		Address = 32'h00000005;
    		#10; 
    		Address = 32'h00000006;
    		#10;
	end
endmodule

